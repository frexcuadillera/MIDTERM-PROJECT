library verilog;
use verilog.vl_types.all;
entity h6to64_tb is
end h6to64_tb;
