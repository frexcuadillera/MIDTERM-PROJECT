library verilog;
use verilog.vl_types.all;
entity binary_encoder83_tb is
end binary_encoder83_tb;
