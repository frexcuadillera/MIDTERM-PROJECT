library verilog;
use verilog.vl_types.all;
entity priority_encoder83_gatelevel_tb is
end priority_encoder83_gatelevel_tb;
