library verilog;
use verilog.vl_types.all;
entity mux41_case_tb is
end mux41_case_tb;
