library verilog;
use verilog.vl_types.all;
entity priority_encoder83_casex_tb is
end priority_encoder83_casex_tb;
