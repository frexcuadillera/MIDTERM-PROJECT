library verilog;
use verilog.vl_types.all;
entity h3to8_tb is
end h3to8_tb;
