//6-to-64 binary decoder
module h6to64(En,w,y);
input En;
input[5:0]w;
input[63:0]y;
wire[7:0]En_w;

h3to8 parent_block(
.En(En),
.w2(w[5]),
.w1(w[4]),
.w0(w[3]),
.y7(En_w[7]),
.y6(En_w[6]),
.y5(En_w[5]),
.y4(En_w[4]),
.y3(En_w[3]),
.y2(En_w[2]),
.y1(En_w[1]),
.y0(En_w[0])
);

h3to8 block0(
.En(En_w[0]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[7]),
.y6(y[6]),
.y5(y[5]),
.y4(y[4]),
.y3(y[3]),
.y2(y[2]),
.y1(y[1]),
.y0(y[0])
);

h3to8 block1(
.En(En_w[1]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[15]),
.y6(y[14]),
.y5(y[13]),
.y4(y[12]),
.y3(y[11]),
.y2(y[10]),
.y1(y[9]),
.y0(y[8])
);

h3to8 block2(
.En(En_w[2]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[23]),
.y6(y[22]),
.y5(y[21]),
.y4(y[20]),
.y3(y[19]),
.y2(y[18]),
.y1(y[17]),
.y0(y[16])
);

h3to8 block3(
.En(En_w[3]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[31]),
.y6(y[30]),
.y5(y[29]),
.y4(y[28]),
.y3(y[27]),
.y2(y[26]),
.y1(y[25]),
.y0(y[24])
);

h3to8 block4(
.En(En_w[4]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[39]),
.y6(y[38]),
.y5(y[37]),
.y4(y[36]),
.y3(y[35]),
.y2(y[34]),
.y1(y[33]),
.y0(y[32])
);

h3to8 block5(
.En(En_w[5]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[47]),
.y6(y[46]),
.y5(y[45]),
.y4(y[44]),
.y3(y[43]),
.y2(y[42]),
.y1(y[41]),
.y0(y[40])
);

h3to8 block6(
.En(En_w[6]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[55]),
.y6(y[54]),
.y5(y[53]),
.y4(y[52]),
.y3(y[51]),
.y2(y[50]),
.y1(y[49]),
.y0(y[48])
);

h3to8 block7(
.En(En_w[7]),
.w2(w[2]),
.w1(w[1]),
.w0(w[0]),
.y7(y[63]),
.y6(y[62]),
.y5(y[61]),
.y4(y[60]),
.y3(y[59]),
.y2(y[58]),
.y1(y[57]),
.y0(y[56])
);
endmodule
