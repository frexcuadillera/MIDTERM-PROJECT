library verilog;
use verilog.vl_types.all;
entity if2to4_tb is
end if2to4_tb;
