library verilog;
use verilog.vl_types.all;
entity binary_encoder42_tb is
end binary_encoder42_tb;
