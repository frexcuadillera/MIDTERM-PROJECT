library verilog;
use verilog.vl_types.all;
entity dec2to4_tb is
end dec2to4_tb;
